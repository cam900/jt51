/*  This file is part of JT51.

    JT51 is free software: you can redistribute it and/or modify
    it under the terms of the GNU General Public License as published by
    the Free Software Foundation, either version 3 of the License, or
    (at your option) any later version.

    JT51 is distributed in the hope that it will be useful,
    but WITHOUT ANY WARRANTY; without even the implied warranty of
    MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
    GNU General Public License for more details.

    You should have received a copy of the GNU General Public License
    along with JT51.  If not, see <http://www.gnu.org/licenses/>.
	
	Author: Jose Tejada Gomez. Twitter: @topapate
	Version: 1.0
	Date: 27-10-2016
	*/
	
10'd0:	 phinc = { 12'd1299	}; // note = 0, KF = 0
10'd1:	 phinc = { 12'd1300	}; // note = 0, KF = 1
10'd2:	 phinc = { 12'd1301	}; // note = 0, KF = 2
10'd3:	 phinc = { 12'd1302	}; // note = 0, KF = 3
10'd4:	 phinc = { 12'd1303	}; // note = 0, KF = 4
10'd5:	 phinc = { 12'd1304	}; // note = 0, KF = 5
10'd6:	 phinc = { 12'd1305	}; // note = 0, KF = 6
10'd7:	 phinc = { 12'd1306	}; // note = 0, KF = 7
10'd8:	 phinc = { 12'd1308	}; // note = 0, KF = 8
10'd9:	 phinc = { 12'd1309	}; // note = 0, KF = 9
10'd10:	 phinc = { 12'd1310	}; // note = 0, KF = 10
10'd11:	 phinc = { 12'd1311	}; // note = 0, KF = 11
10'd12:	 phinc = { 12'd1313	}; // note = 0, KF = 12
10'd13:	 phinc = { 12'd1314	}; // note = 0, KF = 13
10'd14:	 phinc = { 12'd1315	}; // note = 0, KF = 14
10'd15:	 phinc = { 12'd1316	}; // note = 0, KF = 15
10'd16:	 phinc = { 12'd1318	}; // note = 0, KF = 16
10'd17:	 phinc = { 12'd1319	}; // note = 0, KF = 17
10'd18:	 phinc = { 12'd1320	}; // note = 0, KF = 18
10'd19:	 phinc = { 12'd1321	}; // note = 0, KF = 19
10'd20:	 phinc = { 12'd1322	}; // note = 0, KF = 20
10'd21:	 phinc = { 12'd1323	}; // note = 0, KF = 21
10'd22:	 phinc = { 12'd1324	}; // note = 0, KF = 22
10'd23:	 phinc = { 12'd1325	}; // note = 0, KF = 23
10'd24:	 phinc = { 12'd1327	}; // note = 0, KF = 24
10'd25:	 phinc = { 12'd1328	}; // note = 0, KF = 25
10'd26:	 phinc = { 12'd1329	}; // note = 0, KF = 26
10'd27:	 phinc = { 12'd1330	}; // note = 0, KF = 27
10'd28:	 phinc = { 12'd1332	}; // note = 0, KF = 28
10'd29:	 phinc = { 12'd1333	}; // note = 0, KF = 29
10'd30:	 phinc = { 12'd1334	}; // note = 0, KF = 30
10'd31:	 phinc = { 12'd1335	}; // note = 0, KF = 31
10'd32:	 phinc = { 12'd1337	}; // note = 0, KF = 32
10'd33:	 phinc = { 12'd1338	}; // note = 0, KF = 33
10'd34:	 phinc = { 12'd1339	}; // note = 0, KF = 34
10'd35:	 phinc = { 12'd1340	}; // note = 0, KF = 35
10'd36:	 phinc = { 12'd1341	}; // note = 0, KF = 36
10'd37:	 phinc = { 12'd1342	}; // note = 0, KF = 37
10'd38:	 phinc = { 12'd1343	}; // note = 0, KF = 38
10'd39:	 phinc = { 12'd1344	}; // note = 0, KF = 39
10'd40:	 phinc = { 12'd1346	}; // note = 0, KF = 40
10'd41:	 phinc = { 12'd1347	}; // note = 0, KF = 41
10'd42:	 phinc = { 12'd1348	}; // note = 0, KF = 42
10'd43:	 phinc = { 12'd1349	}; // note = 0, KF = 43
10'd44:	 phinc = { 12'd1351	}; // note = 0, KF = 44
10'd45:	 phinc = { 12'd1352	}; // note = 0, KF = 45
10'd46:	 phinc = { 12'd1353	}; // note = 0, KF = 46
10'd47:	 phinc = { 12'd1354	}; // note = 0, KF = 47
10'd48:	 phinc = { 12'd1356	}; // note = 0, KF = 48
10'd49:	 phinc = { 12'd1357	}; // note = 0, KF = 49
10'd50:	 phinc = { 12'd1358	}; // note = 0, KF = 50
10'd51:	 phinc = { 12'd1359	}; // note = 0, KF = 51
10'd52:	 phinc = { 12'd1361	}; // note = 0, KF = 52
10'd53:	 phinc = { 12'd1362	}; // note = 0, KF = 53
10'd54:	 phinc = { 12'd1363	}; // note = 0, KF = 54
10'd55:	 phinc = { 12'd1364	}; // note = 0, KF = 55
10'd56:	 phinc = { 12'd1366	}; // note = 0, KF = 56
10'd57:	 phinc = { 12'd1367	}; // note = 0, KF = 57
10'd58:	 phinc = { 12'd1368	}; // note = 0, KF = 58
10'd59:	 phinc = { 12'd1369	}; // note = 0, KF = 59
10'd60:	 phinc = { 12'd1371	}; // note = 0, KF = 60
10'd61:	 phinc = { 12'd1372	}; // note = 0, KF = 61
10'd62:	 phinc = { 12'd1373	}; // note = 0, KF = 62
10'd63:	 phinc = { 12'd1374	}; // note = 0, KF = 63
10'd64:	 phinc = { 12'd1376	}; // note = 1, KF = 0
10'd65:	 phinc = { 12'd1377	}; // note = 1, KF = 1
10'd66:	 phinc = { 12'd1378	}; // note = 1, KF = 2
10'd67:	 phinc = { 12'd1379	}; // note = 1, KF = 3
10'd68:	 phinc = { 12'd1381	}; // note = 1, KF = 4
10'd69:	 phinc = { 12'd1382	}; // note = 1, KF = 5
10'd70:	 phinc = { 12'd1383	}; // note = 1, KF = 6
10'd71:	 phinc = { 12'd1384	}; // note = 1, KF = 7
10'd72:	 phinc = { 12'd1386	}; // note = 1, KF = 8
10'd73:	 phinc = { 12'd1387	}; // note = 1, KF = 9
10'd74:	 phinc = { 12'd1388	}; // note = 1, KF = 10
10'd75:	 phinc = { 12'd1389	}; // note = 1, KF = 11
10'd76:	 phinc = { 12'd1391	}; // note = 1, KF = 12
10'd77:	 phinc = { 12'd1392	}; // note = 1, KF = 13
10'd78:	 phinc = { 12'd1393	}; // note = 1, KF = 14
10'd79:	 phinc = { 12'd1394	}; // note = 1, KF = 15
10'd80:	 phinc = { 12'd1396	}; // note = 1, KF = 16
10'd81:	 phinc = { 12'd1397	}; // note = 1, KF = 17
10'd82:	 phinc = { 12'd1398	}; // note = 1, KF = 18
10'd83:	 phinc = { 12'd1399	}; // note = 1, KF = 19
10'd84:	 phinc = { 12'd1401	}; // note = 1, KF = 20
10'd85:	 phinc = { 12'd1402	}; // note = 1, KF = 21
10'd86:	 phinc = { 12'd1403	}; // note = 1, KF = 22
10'd87:	 phinc = { 12'd1404	}; // note = 1, KF = 23
10'd88:	 phinc = { 12'd1406	}; // note = 1, KF = 24
10'd89:	 phinc = { 12'd1407	}; // note = 1, KF = 25
10'd90:	 phinc = { 12'd1408	}; // note = 1, KF = 26
10'd91:	 phinc = { 12'd1409	}; // note = 1, KF = 27
10'd92:	 phinc = { 12'd1411	}; // note = 1, KF = 28
10'd93:	 phinc = { 12'd1412	}; // note = 1, KF = 29
10'd94:	 phinc = { 12'd1413	}; // note = 1, KF = 30
10'd95:	 phinc = { 12'd1414	}; // note = 1, KF = 31
10'd96:	 phinc = { 12'd1416	}; // note = 1, KF = 32
10'd97:	 phinc = { 12'd1417	}; // note = 1, KF = 33
10'd98:	 phinc = { 12'd1418	}; // note = 1, KF = 34
10'd99:	 phinc = { 12'd1419	}; // note = 1, KF = 35
10'd100:	 phinc = { 12'd1421	}; // note = 1, KF = 36
10'd101:	 phinc = { 12'd1422	}; // note = 1, KF = 37
10'd102:	 phinc = { 12'd1423	}; // note = 1, KF = 38
10'd103:	 phinc = { 12'd1424	}; // note = 1, KF = 39
10'd104:	 phinc = { 12'd1426	}; // note = 1, KF = 40
10'd105:	 phinc = { 12'd1427	}; // note = 1, KF = 41
10'd106:	 phinc = { 12'd1429	}; // note = 1, KF = 42
10'd107:	 phinc = { 12'd1430	}; // note = 1, KF = 43
10'd108:	 phinc = { 12'd1431	}; // note = 1, KF = 44
10'd109:	 phinc = { 12'd1432	}; // note = 1, KF = 45
10'd110:	 phinc = { 12'd1434	}; // note = 1, KF = 46
10'd111:	 phinc = { 12'd1435	}; // note = 1, KF = 47
10'd112:	 phinc = { 12'd1437	}; // note = 1, KF = 48
10'd113:	 phinc = { 12'd1438	}; // note = 1, KF = 49
10'd114:	 phinc = { 12'd1439	}; // note = 1, KF = 50
10'd115:	 phinc = { 12'd1440	}; // note = 1, KF = 51
10'd116:	 phinc = { 12'd1442	}; // note = 1, KF = 52
10'd117:	 phinc = { 12'd1443	}; // note = 1, KF = 53
10'd118:	 phinc = { 12'd1444	}; // note = 1, KF = 54
10'd119:	 phinc = { 12'd1445	}; // note = 1, KF = 55
10'd120:	 phinc = { 12'd1447	}; // note = 1, KF = 56
10'd121:	 phinc = { 12'd1448	}; // note = 1, KF = 57
10'd122:	 phinc = { 12'd1449	}; // note = 1, KF = 58
10'd123:	 phinc = { 12'd1450	}; // note = 1, KF = 59
10'd124:	 phinc = { 12'd1452	}; // note = 1, KF = 60
10'd125:	 phinc = { 12'd1453	}; // note = 1, KF = 61
10'd126:	 phinc = { 12'd1454	}; // note = 1, KF = 62
10'd127:	 phinc = { 12'd1455	}; // note = 1, KF = 63
10'd128:	 phinc = { 12'd1458	}; // note = 2, KF = 0
10'd129:	 phinc = { 12'd1459	}; // note = 2, KF = 1
10'd130:	 phinc = { 12'd1460	}; // note = 2, KF = 2
10'd131:	 phinc = { 12'd1461	}; // note = 2, KF = 3
10'd132:	 phinc = { 12'd1463	}; // note = 2, KF = 4
10'd133:	 phinc = { 12'd1464	}; // note = 2, KF = 5
10'd134:	 phinc = { 12'd1465	}; // note = 2, KF = 6
10'd135:	 phinc = { 12'd1466	}; // note = 2, KF = 7
10'd136:	 phinc = { 12'd1468	}; // note = 2, KF = 8
10'd137:	 phinc = { 12'd1469	}; // note = 2, KF = 9
10'd138:	 phinc = { 12'd1471	}; // note = 2, KF = 10
10'd139:	 phinc = { 12'd1472	}; // note = 2, KF = 11
10'd140:	 phinc = { 12'd1473	}; // note = 2, KF = 12
10'd141:	 phinc = { 12'd1474	}; // note = 2, KF = 13
10'd142:	 phinc = { 12'd1476	}; // note = 2, KF = 14
10'd143:	 phinc = { 12'd1477	}; // note = 2, KF = 15
10'd144:	 phinc = { 12'd1479	}; // note = 2, KF = 16
10'd145:	 phinc = { 12'd1480	}; // note = 2, KF = 17
10'd146:	 phinc = { 12'd1481	}; // note = 2, KF = 18
10'd147:	 phinc = { 12'd1482	}; // note = 2, KF = 19
10'd148:	 phinc = { 12'd1484	}; // note = 2, KF = 20
10'd149:	 phinc = { 12'd1485	}; // note = 2, KF = 21
10'd150:	 phinc = { 12'd1486	}; // note = 2, KF = 22
10'd151:	 phinc = { 12'd1487	}; // note = 2, KF = 23
10'd152:	 phinc = { 12'd1489	}; // note = 2, KF = 24
10'd153:	 phinc = { 12'd1490	}; // note = 2, KF = 25
10'd154:	 phinc = { 12'd1492	}; // note = 2, KF = 26
10'd155:	 phinc = { 12'd1493	}; // note = 2, KF = 27
10'd156:	 phinc = { 12'd1494	}; // note = 2, KF = 28
10'd157:	 phinc = { 12'd1495	}; // note = 2, KF = 29
10'd158:	 phinc = { 12'd1497	}; // note = 2, KF = 30
10'd159:	 phinc = { 12'd1498	}; // note = 2, KF = 31
10'd160:	 phinc = { 12'd1501	}; // note = 2, KF = 32
10'd161:	 phinc = { 12'd1502	}; // note = 2, KF = 33
10'd162:	 phinc = { 12'd1503	}; // note = 2, KF = 34
10'd163:	 phinc = { 12'd1504	}; // note = 2, KF = 35
10'd164:	 phinc = { 12'd1506	}; // note = 2, KF = 36
10'd165:	 phinc = { 12'd1507	}; // note = 2, KF = 37
10'd166:	 phinc = { 12'd1509	}; // note = 2, KF = 38
10'd167:	 phinc = { 12'd1510	}; // note = 2, KF = 39
10'd168:	 phinc = { 12'd1512	}; // note = 2, KF = 40
10'd169:	 phinc = { 12'd1513	}; // note = 2, KF = 41
10'd170:	 phinc = { 12'd1514	}; // note = 2, KF = 42
10'd171:	 phinc = { 12'd1515	}; // note = 2, KF = 43
10'd172:	 phinc = { 12'd1517	}; // note = 2, KF = 44
10'd173:	 phinc = { 12'd1518	}; // note = 2, KF = 45
10'd174:	 phinc = { 12'd1520	}; // note = 2, KF = 46
10'd175:	 phinc = { 12'd1521	}; // note = 2, KF = 47
10'd176:	 phinc = { 12'd1523	}; // note = 2, KF = 48
10'd177:	 phinc = { 12'd1524	}; // note = 2, KF = 49
10'd178:	 phinc = { 12'd1525	}; // note = 2, KF = 50
10'd179:	 phinc = { 12'd1526	}; // note = 2, KF = 51
10'd180:	 phinc = { 12'd1528	}; // note = 2, KF = 52
10'd181:	 phinc = { 12'd1529	}; // note = 2, KF = 53
10'd182:	 phinc = { 12'd1531	}; // note = 2, KF = 54
10'd183:	 phinc = { 12'd1532	}; // note = 2, KF = 55
10'd184:	 phinc = { 12'd1534	}; // note = 2, KF = 56
10'd185:	 phinc = { 12'd1535	}; // note = 2, KF = 57
10'd186:	 phinc = { 12'd1536	}; // note = 2, KF = 58
10'd187:	 phinc = { 12'd1537	}; // note = 2, KF = 59
10'd188:	 phinc = { 12'd1539	}; // note = 2, KF = 60
10'd189:	 phinc = { 12'd1540	}; // note = 2, KF = 61
10'd190:	 phinc = { 12'd1542	}; // note = 2, KF = 62
10'd191:	 phinc = { 12'd1543	}; // note = 2, KF = 63
10'd192:	 phinc = { 12'd1458	}; // note = 3, KF = 0
10'd193:	 phinc = { 12'd1459	}; // note = 3, KF = 1
10'd194:	 phinc = { 12'd1460	}; // note = 3, KF = 2
10'd195:	 phinc = { 12'd1461	}; // note = 3, KF = 3
10'd196:	 phinc = { 12'd1463	}; // note = 3, KF = 4
10'd197:	 phinc = { 12'd1464	}; // note = 3, KF = 5
10'd198:	 phinc = { 12'd1465	}; // note = 3, KF = 6
10'd199:	 phinc = { 12'd1466	}; // note = 3, KF = 7
10'd200:	 phinc = { 12'd1468	}; // note = 3, KF = 8
10'd201:	 phinc = { 12'd1469	}; // note = 3, KF = 9
10'd202:	 phinc = { 12'd1471	}; // note = 3, KF = 10
10'd203:	 phinc = { 12'd1472	}; // note = 3, KF = 11
10'd204:	 phinc = { 12'd1473	}; // note = 3, KF = 12
10'd205:	 phinc = { 12'd1474	}; // note = 3, KF = 13
10'd206:	 phinc = { 12'd1476	}; // note = 3, KF = 14
10'd207:	 phinc = { 12'd1477	}; // note = 3, KF = 15
10'd208:	 phinc = { 12'd1479	}; // note = 3, KF = 16
10'd209:	 phinc = { 12'd1480	}; // note = 3, KF = 17
10'd210:	 phinc = { 12'd1481	}; // note = 3, KF = 18
10'd211:	 phinc = { 12'd1482	}; // note = 3, KF = 19
10'd212:	 phinc = { 12'd1484	}; // note = 3, KF = 20
10'd213:	 phinc = { 12'd1485	}; // note = 3, KF = 21
10'd214:	 phinc = { 12'd1486	}; // note = 3, KF = 22
10'd215:	 phinc = { 12'd1487	}; // note = 3, KF = 23
10'd216:	 phinc = { 12'd1489	}; // note = 3, KF = 24
10'd217:	 phinc = { 12'd1490	}; // note = 3, KF = 25
10'd218:	 phinc = { 12'd1492	}; // note = 3, KF = 26
10'd219:	 phinc = { 12'd1493	}; // note = 3, KF = 27
10'd220:	 phinc = { 12'd1494	}; // note = 3, KF = 28
10'd221:	 phinc = { 12'd1495	}; // note = 3, KF = 29
10'd222:	 phinc = { 12'd1497	}; // note = 3, KF = 30
10'd223:	 phinc = { 12'd1498	}; // note = 3, KF = 31
10'd224:	 phinc = { 12'd1501	}; // note = 3, KF = 32
10'd225:	 phinc = { 12'd1502	}; // note = 3, KF = 33
10'd226:	 phinc = { 12'd1503	}; // note = 3, KF = 34
10'd227:	 phinc = { 12'd1504	}; // note = 3, KF = 35
10'd228:	 phinc = { 12'd1506	}; // note = 3, KF = 36
10'd229:	 phinc = { 12'd1507	}; // note = 3, KF = 37
10'd230:	 phinc = { 12'd1509	}; // note = 3, KF = 38
10'd231:	 phinc = { 12'd1510	}; // note = 3, KF = 39
10'd232:	 phinc = { 12'd1512	}; // note = 3, KF = 40
10'd233:	 phinc = { 12'd1513	}; // note = 3, KF = 41
10'd234:	 phinc = { 12'd1514	}; // note = 3, KF = 42
10'd235:	 phinc = { 12'd1515	}; // note = 3, KF = 43
10'd236:	 phinc = { 12'd1517	}; // note = 3, KF = 44
10'd237:	 phinc = { 12'd1518	}; // note = 3, KF = 45
10'd238:	 phinc = { 12'd1520	}; // note = 3, KF = 46
10'd239:	 phinc = { 12'd1521	}; // note = 3, KF = 47
10'd240:	 phinc = { 12'd1523	}; // note = 3, KF = 48
10'd241:	 phinc = { 12'd1524	}; // note = 3, KF = 49
10'd242:	 phinc = { 12'd1525	}; // note = 3, KF = 50
10'd243:	 phinc = { 12'd1526	}; // note = 3, KF = 51
10'd244:	 phinc = { 12'd1528	}; // note = 3, KF = 52
10'd245:	 phinc = { 12'd1529	}; // note = 3, KF = 53
10'd246:	 phinc = { 12'd1531	}; // note = 3, KF = 54
10'd247:	 phinc = { 12'd1532	}; // note = 3, KF = 55
10'd248:	 phinc = { 12'd1534	}; // note = 3, KF = 56
10'd249:	 phinc = { 12'd1535	}; // note = 3, KF = 57
10'd250:	 phinc = { 12'd1536	}; // note = 3, KF = 58
10'd251:	 phinc = { 12'd1537	}; // note = 3, KF = 59
10'd252:	 phinc = { 12'd1539	}; // note = 3, KF = 60
10'd253:	 phinc = { 12'd1540	}; // note = 3, KF = 61
10'd254:	 phinc = { 12'd1542	}; // note = 3, KF = 62
10'd255:	 phinc = { 12'd1543	}; // note = 3, KF = 63
10'd256:	 phinc = { 12'd1545	}; // note = 4, KF = 0
10'd257:	 phinc = { 12'd1546	}; // note = 4, KF = 1
10'd258:	 phinc = { 12'd1547	}; // note = 4, KF = 2
10'd259:	 phinc = { 12'd1548	}; // note = 4, KF = 3
10'd260:	 phinc = { 12'd1550	}; // note = 4, KF = 4
10'd261:	 phinc = { 12'd1551	}; // note = 4, KF = 5
10'd262:	 phinc = { 12'd1553	}; // note = 4, KF = 6
10'd263:	 phinc = { 12'd1554	}; // note = 4, KF = 7
10'd264:	 phinc = { 12'd1556	}; // note = 4, KF = 8
10'd265:	 phinc = { 12'd1557	}; // note = 4, KF = 9
10'd266:	 phinc = { 12'd1558	}; // note = 4, KF = 10
10'd267:	 phinc = { 12'd1559	}; // note = 4, KF = 11
10'd268:	 phinc = { 12'd1561	}; // note = 4, KF = 12
10'd269:	 phinc = { 12'd1562	}; // note = 4, KF = 13
10'd270:	 phinc = { 12'd1564	}; // note = 4, KF = 14
10'd271:	 phinc = { 12'd1565	}; // note = 4, KF = 15
10'd272:	 phinc = { 12'd1567	}; // note = 4, KF = 16
10'd273:	 phinc = { 12'd1568	}; // note = 4, KF = 17
10'd274:	 phinc = { 12'd1569	}; // note = 4, KF = 18
10'd275:	 phinc = { 12'd1570	}; // note = 4, KF = 19
10'd276:	 phinc = { 12'd1572	}; // note = 4, KF = 20
10'd277:	 phinc = { 12'd1573	}; // note = 4, KF = 21
10'd278:	 phinc = { 12'd1575	}; // note = 4, KF = 22
10'd279:	 phinc = { 12'd1576	}; // note = 4, KF = 23
10'd280:	 phinc = { 12'd1578	}; // note = 4, KF = 24
10'd281:	 phinc = { 12'd1579	}; // note = 4, KF = 25
10'd282:	 phinc = { 12'd1580	}; // note = 4, KF = 26
10'd283:	 phinc = { 12'd1581	}; // note = 4, KF = 27
10'd284:	 phinc = { 12'd1583	}; // note = 4, KF = 28
10'd285:	 phinc = { 12'd1584	}; // note = 4, KF = 29
10'd286:	 phinc = { 12'd1586	}; // note = 4, KF = 30
10'd287:	 phinc = { 12'd1587	}; // note = 4, KF = 31
10'd288:	 phinc = { 12'd1590	}; // note = 4, KF = 32
10'd289:	 phinc = { 12'd1591	}; // note = 4, KF = 33
10'd290:	 phinc = { 12'd1592	}; // note = 4, KF = 34
10'd291:	 phinc = { 12'd1593	}; // note = 4, KF = 35
10'd292:	 phinc = { 12'd1595	}; // note = 4, KF = 36
10'd293:	 phinc = { 12'd1596	}; // note = 4, KF = 37
10'd294:	 phinc = { 12'd1598	}; // note = 4, KF = 38
10'd295:	 phinc = { 12'd1599	}; // note = 4, KF = 39
10'd296:	 phinc = { 12'd1601	}; // note = 4, KF = 40
10'd297:	 phinc = { 12'd1602	}; // note = 4, KF = 41
10'd298:	 phinc = { 12'd1604	}; // note = 4, KF = 42
10'd299:	 phinc = { 12'd1605	}; // note = 4, KF = 43
10'd300:	 phinc = { 12'd1607	}; // note = 4, KF = 44
10'd301:	 phinc = { 12'd1608	}; // note = 4, KF = 45
10'd302:	 phinc = { 12'd1609	}; // note = 4, KF = 46
10'd303:	 phinc = { 12'd1610	}; // note = 4, KF = 47
10'd304:	 phinc = { 12'd1613	}; // note = 4, KF = 48
10'd305:	 phinc = { 12'd1614	}; // note = 4, KF = 49
10'd306:	 phinc = { 12'd1615	}; // note = 4, KF = 50
10'd307:	 phinc = { 12'd1616	}; // note = 4, KF = 51
10'd308:	 phinc = { 12'd1618	}; // note = 4, KF = 52
10'd309:	 phinc = { 12'd1619	}; // note = 4, KF = 53
10'd310:	 phinc = { 12'd1621	}; // note = 4, KF = 54
10'd311:	 phinc = { 12'd1622	}; // note = 4, KF = 55
10'd312:	 phinc = { 12'd1624	}; // note = 4, KF = 56
10'd313:	 phinc = { 12'd1625	}; // note = 4, KF = 57
10'd314:	 phinc = { 12'd1627	}; // note = 4, KF = 58
10'd315:	 phinc = { 12'd1628	}; // note = 4, KF = 59
10'd316:	 phinc = { 12'd1630	}; // note = 4, KF = 60
10'd317:	 phinc = { 12'd1631	}; // note = 4, KF = 61
10'd318:	 phinc = { 12'd1632	}; // note = 4, KF = 62
10'd319:	 phinc = { 12'd1633	}; // note = 4, KF = 63
10'd320:	 phinc = { 12'd1637	}; // note = 5, KF = 0
10'd321:	 phinc = { 12'd1638	}; // note = 5, KF = 1
10'd322:	 phinc = { 12'd1639	}; // note = 5, KF = 2
10'd323:	 phinc = { 12'd1640	}; // note = 5, KF = 3
10'd324:	 phinc = { 12'd1642	}; // note = 5, KF = 4
10'd325:	 phinc = { 12'd1643	}; // note = 5, KF = 5
10'd326:	 phinc = { 12'd1645	}; // note = 5, KF = 6
10'd327:	 phinc = { 12'd1646	}; // note = 5, KF = 7
10'd328:	 phinc = { 12'd1648	}; // note = 5, KF = 8
10'd329:	 phinc = { 12'd1649	}; // note = 5, KF = 9
10'd330:	 phinc = { 12'd1651	}; // note = 5, KF = 10
10'd331:	 phinc = { 12'd1652	}; // note = 5, KF = 11
10'd332:	 phinc = { 12'd1654	}; // note = 5, KF = 12
10'd333:	 phinc = { 12'd1655	}; // note = 5, KF = 13
10'd334:	 phinc = { 12'd1656	}; // note = 5, KF = 14
10'd335:	 phinc = { 12'd1657	}; // note = 5, KF = 15
10'd336:	 phinc = { 12'd1660	}; // note = 5, KF = 16
10'd337:	 phinc = { 12'd1661	}; // note = 5, KF = 17
10'd338:	 phinc = { 12'd1663	}; // note = 5, KF = 18
10'd339:	 phinc = { 12'd1664	}; // note = 5, KF = 19
10'd340:	 phinc = { 12'd1666	}; // note = 5, KF = 20
10'd341:	 phinc = { 12'd1667	}; // note = 5, KF = 21
10'd342:	 phinc = { 12'd1669	}; // note = 5, KF = 22
10'd343:	 phinc = { 12'd1670	}; // note = 5, KF = 23
10'd344:	 phinc = { 12'd1672	}; // note = 5, KF = 24
10'd345:	 phinc = { 12'd1673	}; // note = 5, KF = 25
10'd346:	 phinc = { 12'd1675	}; // note = 5, KF = 26
10'd347:	 phinc = { 12'd1676	}; // note = 5, KF = 27
10'd348:	 phinc = { 12'd1678	}; // note = 5, KF = 28
10'd349:	 phinc = { 12'd1679	}; // note = 5, KF = 29
10'd350:	 phinc = { 12'd1681	}; // note = 5, KF = 30
10'd351:	 phinc = { 12'd1682	}; // note = 5, KF = 31
10'd352:	 phinc = { 12'd1685	}; // note = 5, KF = 32
10'd353:	 phinc = { 12'd1686	}; // note = 5, KF = 33
10'd354:	 phinc = { 12'd1688	}; // note = 5, KF = 34
10'd355:	 phinc = { 12'd1689	}; // note = 5, KF = 35
10'd356:	 phinc = { 12'd1691	}; // note = 5, KF = 36
10'd357:	 phinc = { 12'd1692	}; // note = 5, KF = 37
10'd358:	 phinc = { 12'd1694	}; // note = 5, KF = 38
10'd359:	 phinc = { 12'd1695	}; // note = 5, KF = 39
10'd360:	 phinc = { 12'd1697	}; // note = 5, KF = 40
10'd361:	 phinc = { 12'd1698	}; // note = 5, KF = 41
10'd362:	 phinc = { 12'd1700	}; // note = 5, KF = 42
10'd363:	 phinc = { 12'd1701	}; // note = 5, KF = 43
10'd364:	 phinc = { 12'd1703	}; // note = 5, KF = 44
10'd365:	 phinc = { 12'd1704	}; // note = 5, KF = 45
10'd366:	 phinc = { 12'd1706	}; // note = 5, KF = 46
10'd367:	 phinc = { 12'd1707	}; // note = 5, KF = 47
10'd368:	 phinc = { 12'd1709	}; // note = 5, KF = 48
10'd369:	 phinc = { 12'd1710	}; // note = 5, KF = 49
10'd370:	 phinc = { 12'd1712	}; // note = 5, KF = 50
10'd371:	 phinc = { 12'd1713	}; // note = 5, KF = 51
10'd372:	 phinc = { 12'd1715	}; // note = 5, KF = 52
10'd373:	 phinc = { 12'd1716	}; // note = 5, KF = 53
10'd374:	 phinc = { 12'd1718	}; // note = 5, KF = 54
10'd375:	 phinc = { 12'd1719	}; // note = 5, KF = 55
10'd376:	 phinc = { 12'd1721	}; // note = 5, KF = 56
10'd377:	 phinc = { 12'd1722	}; // note = 5, KF = 57
10'd378:	 phinc = { 12'd1724	}; // note = 5, KF = 58
10'd379:	 phinc = { 12'd1725	}; // note = 5, KF = 59
10'd380:	 phinc = { 12'd1727	}; // note = 5, KF = 60
10'd381:	 phinc = { 12'd1728	}; // note = 5, KF = 61
10'd382:	 phinc = { 12'd1730	}; // note = 5, KF = 62
10'd383:	 phinc = { 12'd1731	}; // note = 5, KF = 63
10'd384:	 phinc = { 12'd1734	}; // note = 6, KF = 0
10'd385:	 phinc = { 12'd1735	}; // note = 6, KF = 1
10'd386:	 phinc = { 12'd1737	}; // note = 6, KF = 2
10'd387:	 phinc = { 12'd1738	}; // note = 6, KF = 3
10'd388:	 phinc = { 12'd1740	}; // note = 6, KF = 4
10'd389:	 phinc = { 12'd1741	}; // note = 6, KF = 5
10'd390:	 phinc = { 12'd1743	}; // note = 6, KF = 6
10'd391:	 phinc = { 12'd1744	}; // note = 6, KF = 7
10'd392:	 phinc = { 12'd1746	}; // note = 6, KF = 8
10'd393:	 phinc = { 12'd1748	}; // note = 6, KF = 9
10'd394:	 phinc = { 12'd1749	}; // note = 6, KF = 10
10'd395:	 phinc = { 12'd1751	}; // note = 6, KF = 11
10'd396:	 phinc = { 12'd1752	}; // note = 6, KF = 12
10'd397:	 phinc = { 12'd1754	}; // note = 6, KF = 13
10'd398:	 phinc = { 12'd1755	}; // note = 6, KF = 14
10'd399:	 phinc = { 12'd1757	}; // note = 6, KF = 15
10'd400:	 phinc = { 12'd1759	}; // note = 6, KF = 16
10'd401:	 phinc = { 12'd1760	}; // note = 6, KF = 17
10'd402:	 phinc = { 12'd1762	}; // note = 6, KF = 18
10'd403:	 phinc = { 12'd1763	}; // note = 6, KF = 19
10'd404:	 phinc = { 12'd1765	}; // note = 6, KF = 20
10'd405:	 phinc = { 12'd1766	}; // note = 6, KF = 21
10'd406:	 phinc = { 12'd1768	}; // note = 6, KF = 22
10'd407:	 phinc = { 12'd1769	}; // note = 6, KF = 23
10'd408:	 phinc = { 12'd1771	}; // note = 6, KF = 24
10'd409:	 phinc = { 12'd1773	}; // note = 6, KF = 25
10'd410:	 phinc = { 12'd1774	}; // note = 6, KF = 26
10'd411:	 phinc = { 12'd1776	}; // note = 6, KF = 27
10'd412:	 phinc = { 12'd1777	}; // note = 6, KF = 28
10'd413:	 phinc = { 12'd1779	}; // note = 6, KF = 29
10'd414:	 phinc = { 12'd1780	}; // note = 6, KF = 30
10'd415:	 phinc = { 12'd1782	}; // note = 6, KF = 31
10'd416:	 phinc = { 12'd1785	}; // note = 6, KF = 32
10'd417:	 phinc = { 12'd1786	}; // note = 6, KF = 33
10'd418:	 phinc = { 12'd1788	}; // note = 6, KF = 34
10'd419:	 phinc = { 12'd1789	}; // note = 6, KF = 35
10'd420:	 phinc = { 12'd1791	}; // note = 6, KF = 36
10'd421:	 phinc = { 12'd1793	}; // note = 6, KF = 37
10'd422:	 phinc = { 12'd1794	}; // note = 6, KF = 38
10'd423:	 phinc = { 12'd1796	}; // note = 6, KF = 39
10'd424:	 phinc = { 12'd1798	}; // note = 6, KF = 40
10'd425:	 phinc = { 12'd1799	}; // note = 6, KF = 41
10'd426:	 phinc = { 12'd1801	}; // note = 6, KF = 42
10'd427:	 phinc = { 12'd1802	}; // note = 6, KF = 43
10'd428:	 phinc = { 12'd1804	}; // note = 6, KF = 44
10'd429:	 phinc = { 12'd1806	}; // note = 6, KF = 45
10'd430:	 phinc = { 12'd1807	}; // note = 6, KF = 46
10'd431:	 phinc = { 12'd1809	}; // note = 6, KF = 47
10'd432:	 phinc = { 12'd1811	}; // note = 6, KF = 48
10'd433:	 phinc = { 12'd1812	}; // note = 6, KF = 49
10'd434:	 phinc = { 12'd1814	}; // note = 6, KF = 50
10'd435:	 phinc = { 12'd1815	}; // note = 6, KF = 51
10'd436:	 phinc = { 12'd1817	}; // note = 6, KF = 52
10'd437:	 phinc = { 12'd1819	}; // note = 6, KF = 53
10'd438:	 phinc = { 12'd1820	}; // note = 6, KF = 54
10'd439:	 phinc = { 12'd1822	}; // note = 6, KF = 55
10'd440:	 phinc = { 12'd1824	}; // note = 6, KF = 56
10'd441:	 phinc = { 12'd1825	}; // note = 6, KF = 57
10'd442:	 phinc = { 12'd1827	}; // note = 6, KF = 58
10'd443:	 phinc = { 12'd1828	}; // note = 6, KF = 59
10'd444:	 phinc = { 12'd1830	}; // note = 6, KF = 60
10'd445:	 phinc = { 12'd1832	}; // note = 6, KF = 61
10'd446:	 phinc = { 12'd1833	}; // note = 6, KF = 62
10'd447:	 phinc = { 12'd1835	}; // note = 6, KF = 63
10'd448:	 phinc = { 12'd1734	}; // note = 7, KF = 0
10'd449:	 phinc = { 12'd1735	}; // note = 7, KF = 1
10'd450:	 phinc = { 12'd1737	}; // note = 7, KF = 2
10'd451:	 phinc = { 12'd1738	}; // note = 7, KF = 3
10'd452:	 phinc = { 12'd1740	}; // note = 7, KF = 4
10'd453:	 phinc = { 12'd1741	}; // note = 7, KF = 5
10'd454:	 phinc = { 12'd1743	}; // note = 7, KF = 6
10'd455:	 phinc = { 12'd1744	}; // note = 7, KF = 7
10'd456:	 phinc = { 12'd1746	}; // note = 7, KF = 8
10'd457:	 phinc = { 12'd1748	}; // note = 7, KF = 9
10'd458:	 phinc = { 12'd1749	}; // note = 7, KF = 10
10'd459:	 phinc = { 12'd1751	}; // note = 7, KF = 11
10'd460:	 phinc = { 12'd1752	}; // note = 7, KF = 12
10'd461:	 phinc = { 12'd1754	}; // note = 7, KF = 13
10'd462:	 phinc = { 12'd1755	}; // note = 7, KF = 14
10'd463:	 phinc = { 12'd1757	}; // note = 7, KF = 15
10'd464:	 phinc = { 12'd1759	}; // note = 7, KF = 16
10'd465:	 phinc = { 12'd1760	}; // note = 7, KF = 17
10'd466:	 phinc = { 12'd1762	}; // note = 7, KF = 18
10'd467:	 phinc = { 12'd1763	}; // note = 7, KF = 19
10'd468:	 phinc = { 12'd1765	}; // note = 7, KF = 20
10'd469:	 phinc = { 12'd1766	}; // note = 7, KF = 21
10'd470:	 phinc = { 12'd1768	}; // note = 7, KF = 22
10'd471:	 phinc = { 12'd1769	}; // note = 7, KF = 23
10'd472:	 phinc = { 12'd1771	}; // note = 7, KF = 24
10'd473:	 phinc = { 12'd1773	}; // note = 7, KF = 25
10'd474:	 phinc = { 12'd1774	}; // note = 7, KF = 26
10'd475:	 phinc = { 12'd1776	}; // note = 7, KF = 27
10'd476:	 phinc = { 12'd1777	}; // note = 7, KF = 28
10'd477:	 phinc = { 12'd1779	}; // note = 7, KF = 29
10'd478:	 phinc = { 12'd1780	}; // note = 7, KF = 30
10'd479:	 phinc = { 12'd1782	}; // note = 7, KF = 31
10'd480:	 phinc = { 12'd1785	}; // note = 7, KF = 32
10'd481:	 phinc = { 12'd1786	}; // note = 7, KF = 33
10'd482:	 phinc = { 12'd1788	}; // note = 7, KF = 34
10'd483:	 phinc = { 12'd1789	}; // note = 7, KF = 35
10'd484:	 phinc = { 12'd1791	}; // note = 7, KF = 36
10'd485:	 phinc = { 12'd1793	}; // note = 7, KF = 37
10'd486:	 phinc = { 12'd1794	}; // note = 7, KF = 38
10'd487:	 phinc = { 12'd1796	}; // note = 7, KF = 39
10'd488:	 phinc = { 12'd1798	}; // note = 7, KF = 40
10'd489:	 phinc = { 12'd1799	}; // note = 7, KF = 41
10'd490:	 phinc = { 12'd1801	}; // note = 7, KF = 42
10'd491:	 phinc = { 12'd1802	}; // note = 7, KF = 43
10'd492:	 phinc = { 12'd1804	}; // note = 7, KF = 44
10'd493:	 phinc = { 12'd1806	}; // note = 7, KF = 45
10'd494:	 phinc = { 12'd1807	}; // note = 7, KF = 46
10'd495:	 phinc = { 12'd1809	}; // note = 7, KF = 47
10'd496:	 phinc = { 12'd1811	}; // note = 7, KF = 48
10'd497:	 phinc = { 12'd1812	}; // note = 7, KF = 49
10'd498:	 phinc = { 12'd1814	}; // note = 7, KF = 50
10'd499:	 phinc = { 12'd1815	}; // note = 7, KF = 51
10'd500:	 phinc = { 12'd1817	}; // note = 7, KF = 52
10'd501:	 phinc = { 12'd1819	}; // note = 7, KF = 53
10'd502:	 phinc = { 12'd1820	}; // note = 7, KF = 54
10'd503:	 phinc = { 12'd1822	}; // note = 7, KF = 55
10'd504:	 phinc = { 12'd1824	}; // note = 7, KF = 56
10'd505:	 phinc = { 12'd1825	}; // note = 7, KF = 57
10'd506:	 phinc = { 12'd1827	}; // note = 7, KF = 58
10'd507:	 phinc = { 12'd1828	}; // note = 7, KF = 59
10'd508:	 phinc = { 12'd1830	}; // note = 7, KF = 60
10'd509:	 phinc = { 12'd1832	}; // note = 7, KF = 61
10'd510:	 phinc = { 12'd1833	}; // note = 7, KF = 62
10'd511:	 phinc = { 12'd1835	}; // note = 7, KF = 63
10'd512:	 phinc = { 12'd1837	}; // note = 8, KF = 0
10'd513:	 phinc = { 12'd1838	}; // note = 8, KF = 1
10'd514:	 phinc = { 12'd1840	}; // note = 8, KF = 2
10'd515:	 phinc = { 12'd1841	}; // note = 8, KF = 3
10'd516:	 phinc = { 12'd1843	}; // note = 8, KF = 4
10'd517:	 phinc = { 12'd1845	}; // note = 8, KF = 5
10'd518:	 phinc = { 12'd1846	}; // note = 8, KF = 6
10'd519:	 phinc = { 12'd1848	}; // note = 8, KF = 7
10'd520:	 phinc = { 12'd1850	}; // note = 8, KF = 8
10'd521:	 phinc = { 12'd1851	}; // note = 8, KF = 9
10'd522:	 phinc = { 12'd1853	}; // note = 8, KF = 10
10'd523:	 phinc = { 12'd1854	}; // note = 8, KF = 11
10'd524:	 phinc = { 12'd1856	}; // note = 8, KF = 12
10'd525:	 phinc = { 12'd1858	}; // note = 8, KF = 13
10'd526:	 phinc = { 12'd1859	}; // note = 8, KF = 14
10'd527:	 phinc = { 12'd1861	}; // note = 8, KF = 15
10'd528:	 phinc = { 12'd1864	}; // note = 8, KF = 16
10'd529:	 phinc = { 12'd1865	}; // note = 8, KF = 17
10'd530:	 phinc = { 12'd1867	}; // note = 8, KF = 18
10'd531:	 phinc = { 12'd1868	}; // note = 8, KF = 19
10'd532:	 phinc = { 12'd1870	}; // note = 8, KF = 20
10'd533:	 phinc = { 12'd1872	}; // note = 8, KF = 21
10'd534:	 phinc = { 12'd1873	}; // note = 8, KF = 22
10'd535:	 phinc = { 12'd1875	}; // note = 8, KF = 23
10'd536:	 phinc = { 12'd1877	}; // note = 8, KF = 24
10'd537:	 phinc = { 12'd1879	}; // note = 8, KF = 25
10'd538:	 phinc = { 12'd1880	}; // note = 8, KF = 26
10'd539:	 phinc = { 12'd1882	}; // note = 8, KF = 27
10'd540:	 phinc = { 12'd1884	}; // note = 8, KF = 28
10'd541:	 phinc = { 12'd1885	}; // note = 8, KF = 29
10'd542:	 phinc = { 12'd1887	}; // note = 8, KF = 30
10'd543:	 phinc = { 12'd1888	}; // note = 8, KF = 31
10'd544:	 phinc = { 12'd1891	}; // note = 8, KF = 32
10'd545:	 phinc = { 12'd1892	}; // note = 8, KF = 33
10'd546:	 phinc = { 12'd1894	}; // note = 8, KF = 34
10'd547:	 phinc = { 12'd1895	}; // note = 8, KF = 35
10'd548:	 phinc = { 12'd1897	}; // note = 8, KF = 36
10'd549:	 phinc = { 12'd1899	}; // note = 8, KF = 37
10'd550:	 phinc = { 12'd1900	}; // note = 8, KF = 38
10'd551:	 phinc = { 12'd1902	}; // note = 8, KF = 39
10'd552:	 phinc = { 12'd1904	}; // note = 8, KF = 40
10'd553:	 phinc = { 12'd1906	}; // note = 8, KF = 41
10'd554:	 phinc = { 12'd1907	}; // note = 8, KF = 42
10'd555:	 phinc = { 12'd1909	}; // note = 8, KF = 43
10'd556:	 phinc = { 12'd1911	}; // note = 8, KF = 44
10'd557:	 phinc = { 12'd1912	}; // note = 8, KF = 45
10'd558:	 phinc = { 12'd1914	}; // note = 8, KF = 46
10'd559:	 phinc = { 12'd1915	}; // note = 8, KF = 47
10'd560:	 phinc = { 12'd1918	}; // note = 8, KF = 48
10'd561:	 phinc = { 12'd1919	}; // note = 8, KF = 49
10'd562:	 phinc = { 12'd1921	}; // note = 8, KF = 50
10'd563:	 phinc = { 12'd1923	}; // note = 8, KF = 51
10'd564:	 phinc = { 12'd1925	}; // note = 8, KF = 52
10'd565:	 phinc = { 12'd1926	}; // note = 8, KF = 53
10'd566:	 phinc = { 12'd1928	}; // note = 8, KF = 54
10'd567:	 phinc = { 12'd1930	}; // note = 8, KF = 55
10'd568:	 phinc = { 12'd1932	}; // note = 8, KF = 56
10'd569:	 phinc = { 12'd1933	}; // note = 8, KF = 57
10'd570:	 phinc = { 12'd1935	}; // note = 8, KF = 58
10'd571:	 phinc = { 12'd1937	}; // note = 8, KF = 59
10'd572:	 phinc = { 12'd1939	}; // note = 8, KF = 60
10'd573:	 phinc = { 12'd1940	}; // note = 8, KF = 61
10'd574:	 phinc = { 12'd1942	}; // note = 8, KF = 62
10'd575:	 phinc = { 12'd1944	}; // note = 8, KF = 63
10'd576:	 phinc = { 12'd1946	}; // note = 9, KF = 0
10'd577:	 phinc = { 12'd1947	}; // note = 9, KF = 1
10'd578:	 phinc = { 12'd1949	}; // note = 9, KF = 2
10'd579:	 phinc = { 12'd1951	}; // note = 9, KF = 3
10'd580:	 phinc = { 12'd1953	}; // note = 9, KF = 4
10'd581:	 phinc = { 12'd1954	}; // note = 9, KF = 5
10'd582:	 phinc = { 12'd1956	}; // note = 9, KF = 6
10'd583:	 phinc = { 12'd1958	}; // note = 9, KF = 7
10'd584:	 phinc = { 12'd1960	}; // note = 9, KF = 8
10'd585:	 phinc = { 12'd1961	}; // note = 9, KF = 9
10'd586:	 phinc = { 12'd1963	}; // note = 9, KF = 10
10'd587:	 phinc = { 12'd1965	}; // note = 9, KF = 11
10'd588:	 phinc = { 12'd1967	}; // note = 9, KF = 12
10'd589:	 phinc = { 12'd1968	}; // note = 9, KF = 13
10'd590:	 phinc = { 12'd1970	}; // note = 9, KF = 14
10'd591:	 phinc = { 12'd1972	}; // note = 9, KF = 15
10'd592:	 phinc = { 12'd1975	}; // note = 9, KF = 16
10'd593:	 phinc = { 12'd1976	}; // note = 9, KF = 17
10'd594:	 phinc = { 12'd1978	}; // note = 9, KF = 18
10'd595:	 phinc = { 12'd1980	}; // note = 9, KF = 19
10'd596:	 phinc = { 12'd1982	}; // note = 9, KF = 20
10'd597:	 phinc = { 12'd1983	}; // note = 9, KF = 21
10'd598:	 phinc = { 12'd1985	}; // note = 9, KF = 22
10'd599:	 phinc = { 12'd1987	}; // note = 9, KF = 23
10'd600:	 phinc = { 12'd1989	}; // note = 9, KF = 24
10'd601:	 phinc = { 12'd1990	}; // note = 9, KF = 25
10'd602:	 phinc = { 12'd1992	}; // note = 9, KF = 26
10'd603:	 phinc = { 12'd1994	}; // note = 9, KF = 27
10'd604:	 phinc = { 12'd1996	}; // note = 9, KF = 28
10'd605:	 phinc = { 12'd1997	}; // note = 9, KF = 29
10'd606:	 phinc = { 12'd1999	}; // note = 9, KF = 30
10'd607:	 phinc = { 12'd2001	}; // note = 9, KF = 31
10'd608:	 phinc = { 12'd2003	}; // note = 9, KF = 32
10'd609:	 phinc = { 12'd2004	}; // note = 9, KF = 33
10'd610:	 phinc = { 12'd2006	}; // note = 9, KF = 34
10'd611:	 phinc = { 12'd2008	}; // note = 9, KF = 35
10'd612:	 phinc = { 12'd2010	}; // note = 9, KF = 36
10'd613:	 phinc = { 12'd2011	}; // note = 9, KF = 37
10'd614:	 phinc = { 12'd2013	}; // note = 9, KF = 38
10'd615:	 phinc = { 12'd2015	}; // note = 9, KF = 39
10'd616:	 phinc = { 12'd2017	}; // note = 9, KF = 40
10'd617:	 phinc = { 12'd2019	}; // note = 9, KF = 41
10'd618:	 phinc = { 12'd2021	}; // note = 9, KF = 42
10'd619:	 phinc = { 12'd2022	}; // note = 9, KF = 43
10'd620:	 phinc = { 12'd2024	}; // note = 9, KF = 44
10'd621:	 phinc = { 12'd2026	}; // note = 9, KF = 45
10'd622:	 phinc = { 12'd2028	}; // note = 9, KF = 46
10'd623:	 phinc = { 12'd2029	}; // note = 9, KF = 47
10'd624:	 phinc = { 12'd2032	}; // note = 9, KF = 48
10'd625:	 phinc = { 12'd2033	}; // note = 9, KF = 49
10'd626:	 phinc = { 12'd2035	}; // note = 9, KF = 50
10'd627:	 phinc = { 12'd2037	}; // note = 9, KF = 51
10'd628:	 phinc = { 12'd2039	}; // note = 9, KF = 52
10'd629:	 phinc = { 12'd2041	}; // note = 9, KF = 53
10'd630:	 phinc = { 12'd2043	}; // note = 9, KF = 54
10'd631:	 phinc = { 12'd2044	}; // note = 9, KF = 55
10'd632:	 phinc = { 12'd2047	}; // note = 9, KF = 56
10'd633:	 phinc = { 12'd2048	}; // note = 9, KF = 57
10'd634:	 phinc = { 12'd2050	}; // note = 9, KF = 58
10'd635:	 phinc = { 12'd2052	}; // note = 9, KF = 59
10'd636:	 phinc = { 12'd2054	}; // note = 9, KF = 60
10'd637:	 phinc = { 12'd2056	}; // note = 9, KF = 61
10'd638:	 phinc = { 12'd2058	}; // note = 9, KF = 62
10'd639:	 phinc = { 12'd2059	}; // note = 9, KF = 63
10'd640:	 phinc = { 12'd2062	}; // note = 10, KF = 0
10'd641:	 phinc = { 12'd2063	}; // note = 10, KF = 1
10'd642:	 phinc = { 12'd2065	}; // note = 10, KF = 2
10'd643:	 phinc = { 12'd2067	}; // note = 10, KF = 3
10'd644:	 phinc = { 12'd2069	}; // note = 10, KF = 4
10'd645:	 phinc = { 12'd2071	}; // note = 10, KF = 5
10'd646:	 phinc = { 12'd2073	}; // note = 10, KF = 6
10'd647:	 phinc = { 12'd2074	}; // note = 10, KF = 7
10'd648:	 phinc = { 12'd2077	}; // note = 10, KF = 8
10'd649:	 phinc = { 12'd2078	}; // note = 10, KF = 9
10'd650:	 phinc = { 12'd2080	}; // note = 10, KF = 10
10'd651:	 phinc = { 12'd2082	}; // note = 10, KF = 11
10'd652:	 phinc = { 12'd2084	}; // note = 10, KF = 12
10'd653:	 phinc = { 12'd2086	}; // note = 10, KF = 13
10'd654:	 phinc = { 12'd2088	}; // note = 10, KF = 14
10'd655:	 phinc = { 12'd2089	}; // note = 10, KF = 15
10'd656:	 phinc = { 12'd2092	}; // note = 10, KF = 16
10'd657:	 phinc = { 12'd2093	}; // note = 10, KF = 17
10'd658:	 phinc = { 12'd2095	}; // note = 10, KF = 18
10'd659:	 phinc = { 12'd2097	}; // note = 10, KF = 19
10'd660:	 phinc = { 12'd2099	}; // note = 10, KF = 20
10'd661:	 phinc = { 12'd2101	}; // note = 10, KF = 21
10'd662:	 phinc = { 12'd2103	}; // note = 10, KF = 22
10'd663:	 phinc = { 12'd2104	}; // note = 10, KF = 23
10'd664:	 phinc = { 12'd2107	}; // note = 10, KF = 24
10'd665:	 phinc = { 12'd2108	}; // note = 10, KF = 25
10'd666:	 phinc = { 12'd2110	}; // note = 10, KF = 26
10'd667:	 phinc = { 12'd2112	}; // note = 10, KF = 27
10'd668:	 phinc = { 12'd2114	}; // note = 10, KF = 28
10'd669:	 phinc = { 12'd2116	}; // note = 10, KF = 29
10'd670:	 phinc = { 12'd2118	}; // note = 10, KF = 30
10'd671:	 phinc = { 12'd2119	}; // note = 10, KF = 31
10'd672:	 phinc = { 12'd2122	}; // note = 10, KF = 32
10'd673:	 phinc = { 12'd2123	}; // note = 10, KF = 33
10'd674:	 phinc = { 12'd2125	}; // note = 10, KF = 34
10'd675:	 phinc = { 12'd2127	}; // note = 10, KF = 35
10'd676:	 phinc = { 12'd2129	}; // note = 10, KF = 36
10'd677:	 phinc = { 12'd2131	}; // note = 10, KF = 37
10'd678:	 phinc = { 12'd2133	}; // note = 10, KF = 38
10'd679:	 phinc = { 12'd2134	}; // note = 10, KF = 39
10'd680:	 phinc = { 12'd2137	}; // note = 10, KF = 40
10'd681:	 phinc = { 12'd2139	}; // note = 10, KF = 41
10'd682:	 phinc = { 12'd2141	}; // note = 10, KF = 42
10'd683:	 phinc = { 12'd2142	}; // note = 10, KF = 43
10'd684:	 phinc = { 12'd2145	}; // note = 10, KF = 44
10'd685:	 phinc = { 12'd2146	}; // note = 10, KF = 45
10'd686:	 phinc = { 12'd2148	}; // note = 10, KF = 46
10'd687:	 phinc = { 12'd2150	}; // note = 10, KF = 47
10'd688:	 phinc = { 12'd2153	}; // note = 10, KF = 48
10'd689:	 phinc = { 12'd2154	}; // note = 10, KF = 49
10'd690:	 phinc = { 12'd2156	}; // note = 10, KF = 50
10'd691:	 phinc = { 12'd2158	}; // note = 10, KF = 51
10'd692:	 phinc = { 12'd2160	}; // note = 10, KF = 52
10'd693:	 phinc = { 12'd2162	}; // note = 10, KF = 53
10'd694:	 phinc = { 12'd2164	}; // note = 10, KF = 54
10'd695:	 phinc = { 12'd2165	}; // note = 10, KF = 55
10'd696:	 phinc = { 12'd2168	}; // note = 10, KF = 56
10'd697:	 phinc = { 12'd2170	}; // note = 10, KF = 57
10'd698:	 phinc = { 12'd2172	}; // note = 10, KF = 58
10'd699:	 phinc = { 12'd2173	}; // note = 10, KF = 59
10'd700:	 phinc = { 12'd2176	}; // note = 10, KF = 60
10'd701:	 phinc = { 12'd2177	}; // note = 10, KF = 61
10'd702:	 phinc = { 12'd2179	}; // note = 10, KF = 62
10'd703:	 phinc = { 12'd2181	}; // note = 10, KF = 63
10'd704:	 phinc = { 12'd2062	}; // note = 11, KF = 0
10'd705:	 phinc = { 12'd2063	}; // note = 11, KF = 1
10'd706:	 phinc = { 12'd2065	}; // note = 11, KF = 2
10'd707:	 phinc = { 12'd2067	}; // note = 11, KF = 3
10'd708:	 phinc = { 12'd2069	}; // note = 11, KF = 4
10'd709:	 phinc = { 12'd2071	}; // note = 11, KF = 5
10'd710:	 phinc = { 12'd2073	}; // note = 11, KF = 6
10'd711:	 phinc = { 12'd2074	}; // note = 11, KF = 7
10'd712:	 phinc = { 12'd2077	}; // note = 11, KF = 8
10'd713:	 phinc = { 12'd2078	}; // note = 11, KF = 9
10'd714:	 phinc = { 12'd2080	}; // note = 11, KF = 10
10'd715:	 phinc = { 12'd2082	}; // note = 11, KF = 11
10'd716:	 phinc = { 12'd2084	}; // note = 11, KF = 12
10'd717:	 phinc = { 12'd2086	}; // note = 11, KF = 13
10'd718:	 phinc = { 12'd2088	}; // note = 11, KF = 14
10'd719:	 phinc = { 12'd2089	}; // note = 11, KF = 15
10'd720:	 phinc = { 12'd2092	}; // note = 11, KF = 16
10'd721:	 phinc = { 12'd2093	}; // note = 11, KF = 17
10'd722:	 phinc = { 12'd2095	}; // note = 11, KF = 18
10'd723:	 phinc = { 12'd2097	}; // note = 11, KF = 19
10'd724:	 phinc = { 12'd2099	}; // note = 11, KF = 20
10'd725:	 phinc = { 12'd2101	}; // note = 11, KF = 21
10'd726:	 phinc = { 12'd2103	}; // note = 11, KF = 22
10'd727:	 phinc = { 12'd2104	}; // note = 11, KF = 23
10'd728:	 phinc = { 12'd2107	}; // note = 11, KF = 24
10'd729:	 phinc = { 12'd2108	}; // note = 11, KF = 25
10'd730:	 phinc = { 12'd2110	}; // note = 11, KF = 26
10'd731:	 phinc = { 12'd2112	}; // note = 11, KF = 27
10'd732:	 phinc = { 12'd2114	}; // note = 11, KF = 28
10'd733:	 phinc = { 12'd2116	}; // note = 11, KF = 29
10'd734:	 phinc = { 12'd2118	}; // note = 11, KF = 30
10'd735:	 phinc = { 12'd2119	}; // note = 11, KF = 31
10'd736:	 phinc = { 12'd2122	}; // note = 11, KF = 32
10'd737:	 phinc = { 12'd2123	}; // note = 11, KF = 33
10'd738:	 phinc = { 12'd2125	}; // note = 11, KF = 34
10'd739:	 phinc = { 12'd2127	}; // note = 11, KF = 35
10'd740:	 phinc = { 12'd2129	}; // note = 11, KF = 36
10'd741:	 phinc = { 12'd2131	}; // note = 11, KF = 37
10'd742:	 phinc = { 12'd2133	}; // note = 11, KF = 38
10'd743:	 phinc = { 12'd2134	}; // note = 11, KF = 39
10'd744:	 phinc = { 12'd2137	}; // note = 11, KF = 40
10'd745:	 phinc = { 12'd2139	}; // note = 11, KF = 41
10'd746:	 phinc = { 12'd2141	}; // note = 11, KF = 42
10'd747:	 phinc = { 12'd2142	}; // note = 11, KF = 43
10'd748:	 phinc = { 12'd2145	}; // note = 11, KF = 44
10'd749:	 phinc = { 12'd2146	}; // note = 11, KF = 45
10'd750:	 phinc = { 12'd2148	}; // note = 11, KF = 46
10'd751:	 phinc = { 12'd2150	}; // note = 11, KF = 47
10'd752:	 phinc = { 12'd2153	}; // note = 11, KF = 48
10'd753:	 phinc = { 12'd2154	}; // note = 11, KF = 49
10'd754:	 phinc = { 12'd2156	}; // note = 11, KF = 50
10'd755:	 phinc = { 12'd2158	}; // note = 11, KF = 51
10'd756:	 phinc = { 12'd2160	}; // note = 11, KF = 52
10'd757:	 phinc = { 12'd2162	}; // note = 11, KF = 53
10'd758:	 phinc = { 12'd2164	}; // note = 11, KF = 54
10'd759:	 phinc = { 12'd2165	}; // note = 11, KF = 55
10'd760:	 phinc = { 12'd2168	}; // note = 11, KF = 56
10'd761:	 phinc = { 12'd2170	}; // note = 11, KF = 57
10'd762:	 phinc = { 12'd2172	}; // note = 11, KF = 58
10'd763:	 phinc = { 12'd2173	}; // note = 11, KF = 59
10'd764:	 phinc = { 12'd2176	}; // note = 11, KF = 60
10'd765:	 phinc = { 12'd2177	}; // note = 11, KF = 61
10'd766:	 phinc = { 12'd2179	}; // note = 11, KF = 62
10'd767:	 phinc = { 12'd2181	}; // note = 11, KF = 63
10'd768:	 phinc = { 12'd2185	}; // note = 12, KF = 0
10'd769:	 phinc = { 12'd2186	}; // note = 12, KF = 1
10'd770:	 phinc = { 12'd2188	}; // note = 12, KF = 2
10'd771:	 phinc = { 12'd2190	}; // note = 12, KF = 3
10'd772:	 phinc = { 12'd2192	}; // note = 12, KF = 4
10'd773:	 phinc = { 12'd2194	}; // note = 12, KF = 5
10'd774:	 phinc = { 12'd2196	}; // note = 12, KF = 6
10'd775:	 phinc = { 12'd2197	}; // note = 12, KF = 7
10'd776:	 phinc = { 12'd2200	}; // note = 12, KF = 8
10'd777:	 phinc = { 12'd2202	}; // note = 12, KF = 9
10'd778:	 phinc = { 12'd2204	}; // note = 12, KF = 10
10'd779:	 phinc = { 12'd2205	}; // note = 12, KF = 11
10'd780:	 phinc = { 12'd2208	}; // note = 12, KF = 12
10'd781:	 phinc = { 12'd2209	}; // note = 12, KF = 13
10'd782:	 phinc = { 12'd2211	}; // note = 12, KF = 14
10'd783:	 phinc = { 12'd2213	}; // note = 12, KF = 15
10'd784:	 phinc = { 12'd2216	}; // note = 12, KF = 16
10'd785:	 phinc = { 12'd2218	}; // note = 12, KF = 17
10'd786:	 phinc = { 12'd2220	}; // note = 12, KF = 18
10'd787:	 phinc = { 12'd2222	}; // note = 12, KF = 19
10'd788:	 phinc = { 12'd2223	}; // note = 12, KF = 20
10'd789:	 phinc = { 12'd2226	}; // note = 12, KF = 21
10'd790:	 phinc = { 12'd2227	}; // note = 12, KF = 22
10'd791:	 phinc = { 12'd2230	}; // note = 12, KF = 23
10'd792:	 phinc = { 12'd2232	}; // note = 12, KF = 24
10'd793:	 phinc = { 12'd2234	}; // note = 12, KF = 25
10'd794:	 phinc = { 12'd2236	}; // note = 12, KF = 26
10'd795:	 phinc = { 12'd2238	}; // note = 12, KF = 27
10'd796:	 phinc = { 12'd2239	}; // note = 12, KF = 28
10'd797:	 phinc = { 12'd2242	}; // note = 12, KF = 29
10'd798:	 phinc = { 12'd2243	}; // note = 12, KF = 30
10'd799:	 phinc = { 12'd2246	}; // note = 12, KF = 31
10'd800:	 phinc = { 12'd2249	}; // note = 12, KF = 32
10'd801:	 phinc = { 12'd2251	}; // note = 12, KF = 33
10'd802:	 phinc = { 12'd2253	}; // note = 12, KF = 34
10'd803:	 phinc = { 12'd2255	}; // note = 12, KF = 35
10'd804:	 phinc = { 12'd2256	}; // note = 12, KF = 36
10'd805:	 phinc = { 12'd2259	}; // note = 12, KF = 37
10'd806:	 phinc = { 12'd2260	}; // note = 12, KF = 38
10'd807:	 phinc = { 12'd2263	}; // note = 12, KF = 39
10'd808:	 phinc = { 12'd2265	}; // note = 12, KF = 40
10'd809:	 phinc = { 12'd2267	}; // note = 12, KF = 41
10'd810:	 phinc = { 12'd2269	}; // note = 12, KF = 42
10'd811:	 phinc = { 12'd2271	}; // note = 12, KF = 43
10'd812:	 phinc = { 12'd2272	}; // note = 12, KF = 44
10'd813:	 phinc = { 12'd2275	}; // note = 12, KF = 45
10'd814:	 phinc = { 12'd2276	}; // note = 12, KF = 46
10'd815:	 phinc = { 12'd2279	}; // note = 12, KF = 47
10'd816:	 phinc = { 12'd2281	}; // note = 12, KF = 48
10'd817:	 phinc = { 12'd2283	}; // note = 12, KF = 49
10'd818:	 phinc = { 12'd2285	}; // note = 12, KF = 50
10'd819:	 phinc = { 12'd2287	}; // note = 12, KF = 51
10'd820:	 phinc = { 12'd2288	}; // note = 12, KF = 52
10'd821:	 phinc = { 12'd2291	}; // note = 12, KF = 53
10'd822:	 phinc = { 12'd2292	}; // note = 12, KF = 54
10'd823:	 phinc = { 12'd2295	}; // note = 12, KF = 55
10'd824:	 phinc = { 12'd2297	}; // note = 12, KF = 56
10'd825:	 phinc = { 12'd2299	}; // note = 12, KF = 57
10'd826:	 phinc = { 12'd2301	}; // note = 12, KF = 58
10'd827:	 phinc = { 12'd2303	}; // note = 12, KF = 59
10'd828:	 phinc = { 12'd2304	}; // note = 12, KF = 60
10'd829:	 phinc = { 12'd2307	}; // note = 12, KF = 61
10'd830:	 phinc = { 12'd2308	}; // note = 12, KF = 62
10'd831:	 phinc = { 12'd2311	}; // note = 12, KF = 63
10'd832:	 phinc = { 12'd2315	}; // note = 13, KF = 0
10'd833:	 phinc = { 12'd2317	}; // note = 13, KF = 1
10'd834:	 phinc = { 12'd2319	}; // note = 13, KF = 2
10'd835:	 phinc = { 12'd2321	}; // note = 13, KF = 3
10'd836:	 phinc = { 12'd2322	}; // note = 13, KF = 4
10'd837:	 phinc = { 12'd2325	}; // note = 13, KF = 5
10'd838:	 phinc = { 12'd2326	}; // note = 13, KF = 6
10'd839:	 phinc = { 12'd2329	}; // note = 13, KF = 7
10'd840:	 phinc = { 12'd2331	}; // note = 13, KF = 8
10'd841:	 phinc = { 12'd2333	}; // note = 13, KF = 9
10'd842:	 phinc = { 12'd2335	}; // note = 13, KF = 10
10'd843:	 phinc = { 12'd2337	}; // note = 13, KF = 11
10'd844:	 phinc = { 12'd2338	}; // note = 13, KF = 12
10'd845:	 phinc = { 12'd2341	}; // note = 13, KF = 13
10'd846:	 phinc = { 12'd2342	}; // note = 13, KF = 14
10'd847:	 phinc = { 12'd2345	}; // note = 13, KF = 15
10'd848:	 phinc = { 12'd2348	}; // note = 13, KF = 16
10'd849:	 phinc = { 12'd2350	}; // note = 13, KF = 17
10'd850:	 phinc = { 12'd2352	}; // note = 13, KF = 18
10'd851:	 phinc = { 12'd2354	}; // note = 13, KF = 19
10'd852:	 phinc = { 12'd2355	}; // note = 13, KF = 20
10'd853:	 phinc = { 12'd2358	}; // note = 13, KF = 21
10'd854:	 phinc = { 12'd2359	}; // note = 13, KF = 22
10'd855:	 phinc = { 12'd2362	}; // note = 13, KF = 23
10'd856:	 phinc = { 12'd2364	}; // note = 13, KF = 24
10'd857:	 phinc = { 12'd2366	}; // note = 13, KF = 25
10'd858:	 phinc = { 12'd2368	}; // note = 13, KF = 26
10'd859:	 phinc = { 12'd2370	}; // note = 13, KF = 27
10'd860:	 phinc = { 12'd2371	}; // note = 13, KF = 28
10'd861:	 phinc = { 12'd2374	}; // note = 13, KF = 29
10'd862:	 phinc = { 12'd2375	}; // note = 13, KF = 30
10'd863:	 phinc = { 12'd2378	}; // note = 13, KF = 31
10'd864:	 phinc = { 12'd2382	}; // note = 13, KF = 32
10'd865:	 phinc = { 12'd2384	}; // note = 13, KF = 33
10'd866:	 phinc = { 12'd2386	}; // note = 13, KF = 34
10'd867:	 phinc = { 12'd2388	}; // note = 13, KF = 35
10'd868:	 phinc = { 12'd2389	}; // note = 13, KF = 36
10'd869:	 phinc = { 12'd2392	}; // note = 13, KF = 37
10'd870:	 phinc = { 12'd2393	}; // note = 13, KF = 38
10'd871:	 phinc = { 12'd2396	}; // note = 13, KF = 39
10'd872:	 phinc = { 12'd2398	}; // note = 13, KF = 40
10'd873:	 phinc = { 12'd2400	}; // note = 13, KF = 41
10'd874:	 phinc = { 12'd2402	}; // note = 13, KF = 42
10'd875:	 phinc = { 12'd2404	}; // note = 13, KF = 43
10'd876:	 phinc = { 12'd2407	}; // note = 13, KF = 44
10'd877:	 phinc = { 12'd2410	}; // note = 13, KF = 45
10'd878:	 phinc = { 12'd2411	}; // note = 13, KF = 46
10'd879:	 phinc = { 12'd2414	}; // note = 13, KF = 47
10'd880:	 phinc = { 12'd2417	}; // note = 13, KF = 48
10'd881:	 phinc = { 12'd2419	}; // note = 13, KF = 49
10'd882:	 phinc = { 12'd2421	}; // note = 13, KF = 50
10'd883:	 phinc = { 12'd2423	}; // note = 13, KF = 51
10'd884:	 phinc = { 12'd2424	}; // note = 13, KF = 52
10'd885:	 phinc = { 12'd2427	}; // note = 13, KF = 53
10'd886:	 phinc = { 12'd2428	}; // note = 13, KF = 54
10'd887:	 phinc = { 12'd2431	}; // note = 13, KF = 55
10'd888:	 phinc = { 12'd2433	}; // note = 13, KF = 56
10'd889:	 phinc = { 12'd2435	}; // note = 13, KF = 57
10'd890:	 phinc = { 12'd2437	}; // note = 13, KF = 58
10'd891:	 phinc = { 12'd2439	}; // note = 13, KF = 59
10'd892:	 phinc = { 12'd2442	}; // note = 13, KF = 60
10'd893:	 phinc = { 12'd2445	}; // note = 13, KF = 61
10'd894:	 phinc = { 12'd2446	}; // note = 13, KF = 62
10'd895:	 phinc = { 12'd2449	}; // note = 13, KF = 63
10'd896:	 phinc = { 12'd2452	}; // note = 14, KF = 0
10'd897:	 phinc = { 12'd2454	}; // note = 14, KF = 1
10'd898:	 phinc = { 12'd2456	}; // note = 14, KF = 2
10'd899:	 phinc = { 12'd2458	}; // note = 14, KF = 3
10'd900:	 phinc = { 12'd2459	}; // note = 14, KF = 4
10'd901:	 phinc = { 12'd2462	}; // note = 14, KF = 5
10'd902:	 phinc = { 12'd2463	}; // note = 14, KF = 6
10'd903:	 phinc = { 12'd2466	}; // note = 14, KF = 7
10'd904:	 phinc = { 12'd2468	}; // note = 14, KF = 8
10'd905:	 phinc = { 12'd2470	}; // note = 14, KF = 9
10'd906:	 phinc = { 12'd2472	}; // note = 14, KF = 10
10'd907:	 phinc = { 12'd2474	}; // note = 14, KF = 11
10'd908:	 phinc = { 12'd2477	}; // note = 14, KF = 12
10'd909:	 phinc = { 12'd2480	}; // note = 14, KF = 13
10'd910:	 phinc = { 12'd2481	}; // note = 14, KF = 14
10'd911:	 phinc = { 12'd2484	}; // note = 14, KF = 15
10'd912:	 phinc = { 12'd2488	}; // note = 14, KF = 16
10'd913:	 phinc = { 12'd2490	}; // note = 14, KF = 17
10'd914:	 phinc = { 12'd2492	}; // note = 14, KF = 18
10'd915:	 phinc = { 12'd2494	}; // note = 14, KF = 19
10'd916:	 phinc = { 12'd2495	}; // note = 14, KF = 20
10'd917:	 phinc = { 12'd2498	}; // note = 14, KF = 21
10'd918:	 phinc = { 12'd2499	}; // note = 14, KF = 22
10'd919:	 phinc = { 12'd2502	}; // note = 14, KF = 23
10'd920:	 phinc = { 12'd2504	}; // note = 14, KF = 24
10'd921:	 phinc = { 12'd2506	}; // note = 14, KF = 25
10'd922:	 phinc = { 12'd2508	}; // note = 14, KF = 26
10'd923:	 phinc = { 12'd2510	}; // note = 14, KF = 27
10'd924:	 phinc = { 12'd2513	}; // note = 14, KF = 28
10'd925:	 phinc = { 12'd2516	}; // note = 14, KF = 29
10'd926:	 phinc = { 12'd2517	}; // note = 14, KF = 30
10'd927:	 phinc = { 12'd2520	}; // note = 14, KF = 31
10'd928:	 phinc = { 12'd2524	}; // note = 14, KF = 32
10'd929:	 phinc = { 12'd2526	}; // note = 14, KF = 33
10'd930:	 phinc = { 12'd2528	}; // note = 14, KF = 34
10'd931:	 phinc = { 12'd2530	}; // note = 14, KF = 35
10'd932:	 phinc = { 12'd2531	}; // note = 14, KF = 36
10'd933:	 phinc = { 12'd2534	}; // note = 14, KF = 37
10'd934:	 phinc = { 12'd2535	}; // note = 14, KF = 38
10'd935:	 phinc = { 12'd2538	}; // note = 14, KF = 39
10'd936:	 phinc = { 12'd2540	}; // note = 14, KF = 40
10'd937:	 phinc = { 12'd2542	}; // note = 14, KF = 41
10'd938:	 phinc = { 12'd2544	}; // note = 14, KF = 42
10'd939:	 phinc = { 12'd2546	}; // note = 14, KF = 43
10'd940:	 phinc = { 12'd2549	}; // note = 14, KF = 44
10'd941:	 phinc = { 12'd2552	}; // note = 14, KF = 45
10'd942:	 phinc = { 12'd2553	}; // note = 14, KF = 46
10'd943:	 phinc = { 12'd2556	}; // note = 14, KF = 47
10'd944:	 phinc = { 12'd2561	}; // note = 14, KF = 48
10'd945:	 phinc = { 12'd2563	}; // note = 14, KF = 49
10'd946:	 phinc = { 12'd2565	}; // note = 14, KF = 50
10'd947:	 phinc = { 12'd2567	}; // note = 14, KF = 51
10'd948:	 phinc = { 12'd2568	}; // note = 14, KF = 52
10'd949:	 phinc = { 12'd2571	}; // note = 14, KF = 53
10'd950:	 phinc = { 12'd2572	}; // note = 14, KF = 54
10'd951:	 phinc = { 12'd2575	}; // note = 14, KF = 55
10'd952:	 phinc = { 12'd2577	}; // note = 14, KF = 56
10'd953:	 phinc = { 12'd2579	}; // note = 14, KF = 57
10'd954:	 phinc = { 12'd2581	}; // note = 14, KF = 58
10'd955:	 phinc = { 12'd2583	}; // note = 14, KF = 59
10'd956:	 phinc = { 12'd2586	}; // note = 14, KF = 60
10'd957:	 phinc = { 12'd2589	}; // note = 14, KF = 61
10'd958:	 phinc = { 12'd2590	}; // note = 14, KF = 62
10'd959:	 phinc = { 12'd2593	}; // note = 14, KF = 63
10'd960:	 phinc = { 12'd2452	}; // note = 15, KF = 0
10'd961:	 phinc = { 12'd2454	}; // note = 15, KF = 1
10'd962:	 phinc = { 12'd2456	}; // note = 15, KF = 2
10'd963:	 phinc = { 12'd2458	}; // note = 15, KF = 3
10'd964:	 phinc = { 12'd2459	}; // note = 15, KF = 4
10'd965:	 phinc = { 12'd2462	}; // note = 15, KF = 5
10'd966:	 phinc = { 12'd2463	}; // note = 15, KF = 6
10'd967:	 phinc = { 12'd2466	}; // note = 15, KF = 7
10'd968:	 phinc = { 12'd2468	}; // note = 15, KF = 8
10'd969:	 phinc = { 12'd2470	}; // note = 15, KF = 9
10'd970:	 phinc = { 12'd2472	}; // note = 15, KF = 10
10'd971:	 phinc = { 12'd2474	}; // note = 15, KF = 11
10'd972:	 phinc = { 12'd2477	}; // note = 15, KF = 12
10'd973:	 phinc = { 12'd2480	}; // note = 15, KF = 13
10'd974:	 phinc = { 12'd2481	}; // note = 15, KF = 14
10'd975:	 phinc = { 12'd2484	}; // note = 15, KF = 15
10'd976:	 phinc = { 12'd2488	}; // note = 15, KF = 16
10'd977:	 phinc = { 12'd2490	}; // note = 15, KF = 17
10'd978:	 phinc = { 12'd2492	}; // note = 15, KF = 18
10'd979:	 phinc = { 12'd2494	}; // note = 15, KF = 19
10'd980:	 phinc = { 12'd2495	}; // note = 15, KF = 20
10'd981:	 phinc = { 12'd2498	}; // note = 15, KF = 21
10'd982:	 phinc = { 12'd2499	}; // note = 15, KF = 22
10'd983:	 phinc = { 12'd2502	}; // note = 15, KF = 23
10'd984:	 phinc = { 12'd2504	}; // note = 15, KF = 24
10'd985:	 phinc = { 12'd2506	}; // note = 15, KF = 25
10'd986:	 phinc = { 12'd2508	}; // note = 15, KF = 26
10'd987:	 phinc = { 12'd2510	}; // note = 15, KF = 27
10'd988:	 phinc = { 12'd2513	}; // note = 15, KF = 28
10'd989:	 phinc = { 12'd2516	}; // note = 15, KF = 29
10'd990:	 phinc = { 12'd2517	}; // note = 15, KF = 30
10'd991:	 phinc = { 12'd2520	}; // note = 15, KF = 31
10'd992:	 phinc = { 12'd2524	}; // note = 15, KF = 32
10'd993:	 phinc = { 12'd2526	}; // note = 15, KF = 33
10'd994:	 phinc = { 12'd2528	}; // note = 15, KF = 34
10'd995:	 phinc = { 12'd2530	}; // note = 15, KF = 35
10'd996:	 phinc = { 12'd2531	}; // note = 15, KF = 36
10'd997:	 phinc = { 12'd2534	}; // note = 15, KF = 37
10'd998:	 phinc = { 12'd2535	}; // note = 15, KF = 38
10'd999:	 phinc = { 12'd2538	}; // note = 15, KF = 39
10'd1000:	 phinc = { 12'd2540	}; // note = 15, KF = 40
10'd1001:	 phinc = { 12'd2542	}; // note = 15, KF = 41
10'd1002:	 phinc = { 12'd2544	}; // note = 15, KF = 42
10'd1003:	 phinc = { 12'd2546	}; // note = 15, KF = 43
10'd1004:	 phinc = { 12'd2549	}; // note = 15, KF = 44
10'd1005:	 phinc = { 12'd2552	}; // note = 15, KF = 45
10'd1006:	 phinc = { 12'd2553	}; // note = 15, KF = 46
10'd1007:	 phinc = { 12'd2556	}; // note = 15, KF = 47
10'd1008:	 phinc = { 12'd2561	}; // note = 15, KF = 48
10'd1009:	 phinc = { 12'd2563	}; // note = 15, KF = 49
10'd1010:	 phinc = { 12'd2565	}; // note = 15, KF = 50
10'd1011:	 phinc = { 12'd2567	}; // note = 15, KF = 51
10'd1012:	 phinc = { 12'd2568	}; // note = 15, KF = 52
10'd1013:	 phinc = { 12'd2571	}; // note = 15, KF = 53
10'd1014:	 phinc = { 12'd2572	}; // note = 15, KF = 54
10'd1015:	 phinc = { 12'd2575	}; // note = 15, KF = 55
10'd1016:	 phinc = { 12'd2577	}; // note = 15, KF = 56
10'd1017:	 phinc = { 12'd2579	}; // note = 15, KF = 57
10'd1018:	 phinc = { 12'd2581	}; // note = 15, KF = 58
10'd1019:	 phinc = { 12'd2583	}; // note = 15, KF = 59
10'd1020:	 phinc = { 12'd2586	}; // note = 15, KF = 60
10'd1021:	 phinc = { 12'd2589	}; // note = 15, KF = 61
10'd1022:	 phinc = { 12'd2590	}; // note = 15, KF = 62
10'd1023:	 phinc = { 12'd2593	}; // note = 15, KF = 63
